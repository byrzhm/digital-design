module my_design;

    task print;
        $display("I'm at %m");
    endtask

endmodule
